//7 segments digits

`define ZERO    8'b10001000
`define ONE     8'b11111001
`define TWO     8'b01001100
`define THREE   8'b01101000
`define FOUR    8'b10011001
`define FIVE    8'b00101010
`define SIX     8'b00001010
`define SEVEN   8'b11111000
`define EIGHT   8'b00001000
`define NINE    8'b00101000
