module hello;
  initial
    begin
      $display("Hello Mario");
      $finish ;
    end
endmodule
