`default_nettype none

module rom32x4 (input clk,
				input wire [4:0] addr,
				output reg [3:0]data);

	reg [3:0] rom [0:31];

	always @(negedge clk) begin
		data <= rom[addr];
	end

	initial begin
		rom[0] = 4'h0; 
	    rom[1] = 4'h1;
	    rom[2] = 4'h2;
	    rom[3] = 4'h3;
	    rom[4] = 4'h4; 
	    rom[5] = 4'h5;
	    rom[6] = 4'h6;
	    rom[7] = 4'h7;
	end

endmodule